-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION vm_circuit_beta_struct_config OF vm_circuit_beta IS
   FOR struct
   END FOR;
END vm_circuit_beta_struct_config;
