-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION next_state_logic_struct_config OF next_state_logic IS
   FOR struct
   END FOR;
END next_state_logic_struct_config;
