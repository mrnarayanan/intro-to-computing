-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION nextstatelogic_beta_struct_config OF nextstatelogic_beta IS
   FOR struct
   END FOR;
END nextstatelogic_beta_struct_config;
